VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END Y
END AND2x2

MACRO AND3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.344 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END Y
END AND3x1

MACRO AND3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2 0 0 ;
SIZE 1.512 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END Y
END AND3x2

MACRO AOI21x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1 0 0 ;
SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.52 0.576 0.776 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.52 0.144 0.776 ;
    END
  END Y
END AOI21x1

MACRO AOI22x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22x1 0 0 ;
SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.52 0.36 0.776 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.344 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.52 0.576 0.776 ;
    END
  END Y
END AOI22x1

MACRO BUFx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2 0 0 ;
SIZE 1.08 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END Y
END BUFx2

MACRO BUFx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END Y
END BUFx3

MACRO BUFx4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4 0 0 ;
SIZE 1.512 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END Y
END BUFx4

MACRO BUFx8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8 0 0 ;
SIZE 2.592 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.232 0.088 2.304 0.344 ;
    END
  END Y
END BUFx8

MACRO DFFHQNx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx1 0 0 ;
SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 0.072 0.52 0.144 0.776 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.344 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.088 1.656 0.344 ;
    END
  END QN
  OBS
    LAYER M1 ;
RECT 1.8 0.232 1.872 0.776 ;
RECT 1.584 0.52 1.656 0.776 ;
RECT 1.368 0.088 1.44 0.776 ;
RECT 1.152 0.232 1.224 0.632 ;
RECT 0.936 0.52 1.008 0.776 ;
RECT 0.72 0.088 0.792 0.344 ;
RECT 0.72 0.52 0.792 0.776 ;
RECT 0.504 0.52 0.576 0.776 ;
RECT 0.288 0.232 0.36 0.632 ;
    LAYER M2 ;
RECT 0.916 0.54 1.892 0.612 ;
RECT 0.484 0.684 1.676 0.756 ;
    LAYER V1 ;
RECT 1.8 0.54 1.872 0.612 ;
RECT 1.584 0.684 1.656 0.756 ;
RECT 0.936 0.54 1.008 0.612 ;
RECT 0.504 0.684 0.576 0.756 ;
  END
END DFFHQNx1

MACRO DFFHQNx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx2 0 0 ;
SIZE 1.944 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 1.584 0.52 1.656 0.776 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.52 1.008 0.776 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.52 1.224 0.776 ;
    END
  END QN
  OBS
    LAYER M1 ;
RECT 1.8 0.088 1.872 0.632 ;
RECT 1.584 0.088 1.656 0.344 ;
RECT 1.368 0.232 1.44 0.776 ;
RECT 0.72 0.088 0.792 0.776 ;
RECT 0.288 0.232 0.36 0.632 ;
RECT 0.072 0.088 0.144 0.776 ;
    LAYER M2 ;
RECT 0.7 0.108 1.676 0.18 ;
    LAYER V1 ;
RECT 1.584 0.108 1.656 0.18 ;
RECT 0.72 0.108 0.792 0.18 ;
  END
END DFFHQNx2

MACRO DFFHQNx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx3 0 0 ;
SIZE 2.16 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 1.584 0.52 1.656 0.776 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
    END
  END QN
  OBS
    LAYER M1 ;
RECT 2.016 0.088 2.088 0.632 ;
RECT 1.8 0.232 1.872 0.776 ;
RECT 1.584 0.088 1.656 0.344 ;
RECT 1.368 0.232 1.44 0.776 ;
RECT 0.72 0.088 0.792 0.776 ;
RECT 0.504 0.232 0.576 0.632 ;
RECT 0.288 0.232 0.36 0.776 ;
RECT 0.072 0.088 0.144 0.632 ;
    LAYER M2 ;
RECT 0.484 0.252 1.892 0.324 ;
    LAYER V1 ;
RECT 1.8 0.252 1.872 0.324 ;
RECT 1.584 0.252 1.656 0.324 ;
RECT 0.504 0.252 0.576 0.324 ;
  END
END DFFHQNx3

MACRO DHLx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx1 0 0 ;
SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.52 0.144 0.776 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END Q
  OBS
    LAYER M1 ;
RECT 1.368 0.232 1.44 0.632 ;
RECT 0.936 0.232 1.008 0.632 ;
RECT 0.72 0.232 0.792 0.632 ;
RECT 0.504 0.088 0.576 0.776 ;
RECT 0.288 0.232 0.36 0.632 ;
    LAYER M2 ;
RECT 0.268 0.252 1.028 0.324 ;
    LAYER V1 ;
RECT 0.936 0.252 1.008 0.324 ;
RECT 0.288 0.252 0.36 0.324 ;
  END
END DHLx1

MACRO DHLx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx2 0 0 ;
SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 1.152 0.52 1.224 0.776 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.52 0.36 0.776 ;
    END
  END Q
  OBS
    LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
RECT 0.936 0.232 1.008 0.632 ;
RECT 0.72 0.088 0.792 0.776 ;
RECT 0.504 0.232 0.576 0.632 ;
RECT 0.072 0.232 0.144 0.632 ;
    LAYER M2 ;
RECT 0.052 0.252 1.244 0.324 ;
    LAYER V1 ;
RECT 1.152 0.252 1.224 0.324 ;
RECT 0.072 0.252 0.144 0.324 ;
  END
END DHLx2

MACRO DHLx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx3 0 0 ;
SIZE 1.728 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 0.936 0.52 1.008 0.776 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.088 1.44 0.344 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END Q
  OBS
    LAYER M1 ;
RECT 1.152 0.088 1.224 0.632 ;
RECT 0.936 0.088 1.008 0.344 ;
RECT 0.72 0.232 0.792 0.632 ;
RECT 0.504 0.232 0.576 0.776 ;
    LAYER M2 ;
RECT 0.7 0.252 1.028 0.324 ;
    LAYER V1 ;
RECT 0.936 0.252 1.008 0.324 ;
RECT 0.72 0.252 0.792 0.324 ;
  END
END DHLx3

MACRO FAx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FAx1 0 0 ;
SIZE 1.512 BY 1.296 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.52 1.224 1.064 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 1.064 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 1.064 ;
    END
  END CI
  PIN CON
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.232 1.44 1.064 ;
    END
  END CON
  PIN SN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.952 0.144 1.208 ;
    END
  END SN
  OBS
    LAYER M1 ;
RECT 0.936 0.232 1.008 0.776 ;
  END
END FAx1

MACRO INVx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1 0 0 ;
SIZE 0.648 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END Y
END INVx1

MACRO INVx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2 0 0 ;
SIZE 0.864 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.344 ;
    END
  END Y
END INVx2

MACRO INVx4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END Y
END INVx4

MACRO INVx8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8 0 0 ;
SIZE 2.16 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.088 1.872 0.344 ;
    END
  END Y
END INVx8

MACRO NAND2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
RECT 0.484 0.252 1.244 0.324 ;
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
RECT 0.504 0.088 0.576 0.344 ;
      LAYER V1 ;
RECT 0.504 0.252 0.576 0.324 ;
RECT 1.152 0.252 1.224 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
RECT 0.288 0.088 0.36 0.344 ;
    LAYER M2 ;
RECT 0.268 0.108 0.812 0.18 ;
    LAYER V1 ;
RECT 0.72 0.108 0.792 0.18 ;
RECT 0.288 0.108 0.36 0.18 ;
  END
END NAND2x1

MACRO NAND2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2 0 0 ;
SIZE 2.16 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.088 1.872 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
RECT 0.484 0.108 1.46 0.18 ;
      LAYER M1 ;
RECT 1.368 0.088 1.44 0.344 ;
RECT 0.936 0.088 1.008 0.344 ;
RECT 0.504 0.088 0.576 0.344 ;
      LAYER V1 ;
RECT 0.504 0.108 0.576 0.18 ;
RECT 0.936 0.108 1.008 0.18 ;
RECT 1.368 0.108 1.44 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 1.584 0.088 1.656 0.344 ;
RECT 1.152 0.088 1.224 0.344 ;
RECT 0.72 0.088 0.792 0.344 ;
RECT 0.288 0.088 0.36 0.344 ;
    LAYER M2 ;
RECT 0.268 0.252 1.676 0.324 ;
    LAYER V1 ;
RECT 1.584 0.252 1.656 0.324 ;
RECT 1.152 0.252 1.224 0.324 ;
RECT 0.72 0.252 0.792 0.324 ;
RECT 0.288 0.252 0.36 0.324 ;
  END
END NAND2x2

MACRO NAND3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1 0 0 ;
SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.52 1.224 0.776 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.52 0.792 0.776 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
RECT 0.484 0.252 1.244 0.324 ;
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
RECT 0.936 0.088 1.008 0.344 ;
RECT 0.504 0.088 0.576 0.344 ;
      LAYER V1 ;
RECT 0.504 0.252 0.576 0.324 ;
RECT 0.936 0.252 1.008 0.324 ;
RECT 1.152 0.252 1.224 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
RECT 0.288 0.088 0.36 0.344 ;
    LAYER M2 ;
RECT 0.268 0.108 0.812 0.18 ;
    LAYER V1 ;
RECT 0.72 0.108 0.792 0.18 ;
RECT 0.288 0.108 0.36 0.18 ;
  END
END NAND3x1

MACRO NAND3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2 0 0 ;
SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.52 0.36 0.776 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.52 1.008 0.776 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.52 1.656 0.776 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.016 0.232 2.088 0.632 ;
    END
  END Y
END NAND3x2

MACRO NOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
RECT 0.052 0.108 0.812 0.18 ;
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
RECT 0.072 0.088 0.144 0.344 ;
      LAYER V1 ;
RECT 0.072 0.108 0.144 0.18 ;
RECT 0.72 0.108 0.792 0.18 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
RECT 0.504 0.088 0.576 0.344 ;
    LAYER M2 ;
RECT 0.484 0.252 1.244 0.324 ;
    LAYER V1 ;
RECT 1.152 0.252 1.224 0.324 ;
RECT 0.504 0.252 0.576 0.324 ;
  END
END NOR2x1

MACRO NOR2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2 0 0 ;
SIZE 2.16 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.088 1.872 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
RECT 0.484 0.252 1.676 0.324 ;
      LAYER M1 ;
RECT 1.584 0.088 1.656 0.344 ;
RECT 1.152 0.088 1.224 0.344 ;
RECT 0.504 0.088 0.576 0.344 ;
      LAYER V1 ;
RECT 0.504 0.252 0.576 0.324 ;
RECT 1.152 0.252 1.224 0.324 ;
RECT 1.584 0.252 1.656 0.324 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 2.016 0.088 2.088 0.344 ;
RECT 1.368 0.088 1.44 0.344 ;
RECT 0.936 0.088 1.008 0.344 ;
RECT 0.72 0.088 0.792 0.344 ;
RECT 0.288 0.088 0.36 0.344 ;
    LAYER M2 ;
RECT 0.916 0.108 2.108 0.18 ;
RECT 0.268 0.108 0.812 0.18 ;
    LAYER V1 ;
RECT 2.016 0.108 2.088 0.18 ;
RECT 1.368 0.108 1.44 0.18 ;
RECT 0.936 0.108 1.008 0.18 ;
RECT 0.72 0.108 0.792 0.18 ;
RECT 0.288 0.108 0.36 0.18 ;
  END
END NOR2x2

MACRO NOR3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1 0 0 ;
SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.52 0.144 0.776 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
RECT 0.484 0.684 1.244 0.756 ;
      LAYER M1 ;
RECT 1.152 0.52 1.224 0.776 ;
RECT 0.936 0.52 1.008 0.776 ;
RECT 0.504 0.52 0.576 0.776 ;
      LAYER V1 ;
RECT 0.504 0.684 0.576 0.756 ;
RECT 0.936 0.684 1.008 0.756 ;
RECT 1.152 0.684 1.224 0.756 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 0.72 0.52 0.792 0.776 ;
RECT 0.288 0.232 0.36 0.632 ;
    LAYER M2 ;
RECT 0.268 0.54 0.812 0.612 ;
    LAYER V1 ;
RECT 0.72 0.54 0.792 0.612 ;
RECT 0.288 0.54 0.36 0.612 ;
  END
END NOR3x1

MACRO NOR3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2 0 0 ;
SIZE 2.376 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.016 0.088 2.088 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.776 ;
    END
  END Y
END NOR3x2

MACRO OAI21x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21x1 0 0 ;
SIZE 1.08 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.52 0.792 0.776 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 0.632 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.52 0.36 0.776 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
  END
END OAI21x1

MACRO OAI22x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22x1 0 0 ;
SIZE 1.296 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.52 0.36 0.776 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.344 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.52 0.792 0.776 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 0.504 0.52 0.576 0.776 ;
  END
END OAI22x1

MACRO OR2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END Y
END OR2x2

MACRO OR3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1 0 0 ;
SIZE 1.296 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.344 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.344 ;
    END
  END Y
END OR3x1

MACRO OR3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2 0 0 ;
SIZE 1.512 BY 0.432 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.344 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.344 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END Y
END OR3x2

MACRO XNOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x1 0 0 ;
SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.344 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.52 0.576 0.776 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.344 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 0.936 0.232 1.008 0.776 ;
RECT 0.288 0.52 0.36 0.776 ;
  END
END XNOR2x1

MACRO XOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x1 0 0 ;
SIZE 1.512 BY 0.864 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.52 0.36 0.776 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.232 1.224 0.632 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
RECT 0.484 0.252 0.812 0.324 ;
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
RECT 0.504 0.088 0.576 0.344 ;
      LAYER V1 ;
RECT 0.504 0.252 0.576 0.324 ;
RECT 0.72 0.252 0.792 0.324 ;
    END
  END Y
END XOR2x1

END LIBRARY
