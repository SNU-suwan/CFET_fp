VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.488 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 0.632 ;
    END
  END Y
END AND2x2

MACRO AND3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.488 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 0.632 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END Y
END AND3x1

MACRO AND3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2 0 0 ;
SIZE 1.512 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.232 1.224 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.488 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END Y
END AND3x2

MACRO AOI21x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1 0 0 ;
SIZE 1.944 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.088 1.44 0.488 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.488 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END Y
END AOI21x1

MACRO AOI22x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22x1 0 0 ;
SIZE 2.376 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.232 1.44 0.632 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.016 0.088 2.088 0.488 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.488 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 1.8 0.376 1.872 0.632 ;
RECT 0.504 0.376 0.576 0.632 ;
    LAYER M2 ;
RECT 0.484 0.54 1.892 0.612 ;
    LAYER V1 ;
RECT 1.8 0.54 1.872 0.612 ;
RECT 0.504 0.54 0.576 0.612 ;
  END
END AOI22x1

MACRO BUFx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2 0 0 ;
SIZE 1.08 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END Y
END BUFx2

MACRO BUFx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END Y
END BUFx3

MACRO BUFx4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4 0 0 ;
SIZE 1.512 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.488 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 0.632 ;
    END
  END Y
END BUFx4

MACRO BUFx8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8 0 0 ;
SIZE 2.592 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.232 1.872 0.632 ;
    END
  END Y
END BUFx8

MACRO DFFHQNx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx1 0 0 ;
SIZE 3.24 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.488 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END QN
  OBS
    LAYER M1 ;
RECT 2.232 0.232 2.304 0.488 ;
RECT 1.584 0.232 1.656 0.488 ;
    LAYER M2 ;
RECT 1.564 0.252 2.324 0.324 ;
    LAYER V1 ;
RECT 2.232 0.252 2.304 0.324 ;
RECT 1.584 0.252 1.656 0.324 ;
  END
END DFFHQNx1

MACRO DFFHQNx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx2 0 0 ;
SIZE 3.456 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 3.096 0.232 3.168 0.632 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.232 0.232 2.304 0.632 ;
    END
  END QN
  OBS
    LAYER M1 ;
RECT 2.448 0.376 2.52 0.632 ;
RECT 1.8 0.376 1.872 0.632 ;
    LAYER M2 ;
RECT 1.78 0.396 2.54 0.468 ;
    LAYER V1 ;
RECT 2.448 0.396 2.52 0.468 ;
RECT 1.8 0.396 1.872 0.468 ;
  END
END DFFHQNx2

MACRO DFFHQNx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx3 0 0 ;
SIZE 3.672 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.088 1.656 0.488 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END QN
  OBS
    LAYER M1 ;
RECT 2.664 0.232 2.736 0.488 ;
RECT 2.016 0.088 2.088 0.344 ;
    LAYER M2 ;
RECT 1.996 0.252 2.756 0.324 ;
    LAYER V1 ;
RECT 2.664 0.252 2.736 0.324 ;
RECT 2.016 0.252 2.088 0.324 ;
  END
END DFFHQNx3

MACRO DHLx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx1 0 0 ;
SIZE 2.376 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.088 1.872 0.488 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.016 0.232 2.088 0.632 ;
    END
  END Q
END DHLx1

MACRO DHLx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx2 0 0 ;
SIZE 2.592 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.232 1.872 0.632 ;
    END
  END Q
END DHLx2

MACRO DHLx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx3 0 0 ;
SIZE 2.808 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION OUTPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
RECT 1.368 0.232 1.44 0.632 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.232 0.088 2.304 0.488 ;
    END
  END D
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END Q
END DHLx3

MACRO INVx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1 0 0 ;
SIZE 0.648 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.232 0.144 0.632 ;
    END
  END Y
END INVx1

MACRO INVx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2 0 0 ;
SIZE 0.864 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 0.632 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END Y
END INVx2

MACRO INVx4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.488 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END Y
END INVx4

MACRO INVx8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8 0 0 ;
SIZE 2.16 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.232 0.144 0.632 ;
    END
  END Y
END INVx8

MACRO NAND2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.488 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 0.632 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END Y
END NAND2x1

MACRO NAND2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2 0 0 ;
SIZE 2.16 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.232 1.872 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END Y
END NAND2x2

MACRO NAND3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1 0 0 ;
SIZE 2.376 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.232 1.44 0.632 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.232 1.656 0.632 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.016 0.088 2.088 0.488 ;
    END
  END Y
END NAND3x1

MACRO NAND3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2 0 0 ;
SIZE 4.536 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.088 1.44 0.488 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 3.096 0.088 3.168 0.488 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.88 0.088 2.952 0.488 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.232 0.144 0.632 ;
    END
  END Y
END NAND3x2

MACRO NOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.488 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.488 ;
    END
  END Y
END NOR2x1

MACRO NOR2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2 0 0 ;
SIZE 2.16 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.088 0.36 0.488 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.088 1.224 0.488 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.232 1.872 0.632 ;
    END
  END Y
END NOR2x2

MACRO NOR3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1 0 0 ;
SIZE 2.376 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 2.016 0.232 2.088 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 1.8 0.088 1.872 0.632 ;
  END
END NOR3x1

MACRO NOR3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2 0 0 ;
SIZE 4.536 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.232 1.872 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 4.176 0.232 4.248 0.632 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.232 1.44 0.632 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.488 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 2.88 0.232 2.952 0.632 ;
RECT 2.664 0.088 2.736 0.632 ;
RECT 2.448 0.088 2.52 0.344 ;
    LAYER M2 ;
RECT 2.428 0.252 2.972 0.324 ;
    LAYER V1 ;
RECT 2.88 0.252 2.952 0.324 ;
RECT 2.448 0.252 2.52 0.324 ;
  END
END NOR3x2

MACRO OAI21x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21x1 0 0 ;
SIZE 1.944 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.488 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.088 1.44 0.488 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.232 1.656 0.632 ;
    END
  END Y
END OAI21x1

MACRO OAI22x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22x1 0 0 ;
SIZE 2.376 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.232 0.576 0.632 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.8 0.088 1.872 0.488 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.368 0.232 1.44 0.632 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.088 1.656 0.488 ;
    END
  END Y
END OAI22x1

MACRO OR2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.088 1.008 0.488 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END Y
END OR2x2

MACRO OR3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1 0 0 ;
SIZE 1.296 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.488 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.504 0.088 0.576 0.488 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.488 ;
    END
  END Y
END OR3x1

MACRO OR3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2 0 0 ;
SIZE 1.512 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.152 0.232 1.224 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.936 0.232 1.008 0.632 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.088 0.792 0.488 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END Y
END OR3x2

MACRO XNOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x1 0 0 ;
SIZE 2.376 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.232 1.656 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.288 0.232 0.36 0.632 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.088 0.144 0.488 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 1.368 0.088 1.44 0.488 ;
RECT 0.504 0.376 0.576 0.632 ;
    LAYER M2 ;
RECT 0.484 0.396 1.46 0.468 ;
    LAYER V1 ;
RECT 1.368 0.396 1.44 0.468 ;
RECT 0.504 0.396 0.576 0.468 ;
  END
END XNOR2x1

MACRO XOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x1 0 0 ;
SIZE 2.376 BY 0.72 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 1.584 0.232 1.656 0.632 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.72 0.232 0.792 0.632 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
RECT 0.072 0.232 0.144 0.632 ;
    END
  END Y
  OBS
    LAYER M1 ;
RECT 1.368 0.376 1.44 0.632 ;
RECT 0.504 0.232 0.576 0.488 ;
    LAYER M2 ;
RECT 0.484 0.396 1.46 0.468 ;
    LAYER V1 ;
RECT 1.368 0.396 1.44 0.468 ;
RECT 0.504 0.396 0.576 0.468 ;
  END
END XOR2x1

END LIBRARY
