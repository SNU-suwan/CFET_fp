VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Y
END AND2x2

MACRO AND3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END Y
END AND3x1

MACRO AND3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2 0 0 ;
  SIZE 0.378 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END Y
END AND3x2

MACRO AOI21x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1 0 0 ;
  SIZE 0.486 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.022 0.36 0.122 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.175 0.099 0.311 0.117 ;
      LAYER M1 ;
        RECT 0.288 0.058 0.306 0.122 ;
        RECT 0.18 0.022 0.198 0.122 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
        RECT 0.288 0.099 0.306 0.117 ;
    END
  END Y
END AOI21x1

MACRO AOI22x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22x1 0 0 ;
  SIZE 0.648 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.022 0.522 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.022 0.414 0.122 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.121 0.099 0.365 0.117 ;
      LAYER M1 ;
        RECT 0.342 0.058 0.36 0.122 ;
        RECT 0.126 0.022 0.144 0.122 ;
      LAYER V1 ;
        RECT 0.126 0.099 0.144 0.117 ;
        RECT 0.342 0.099 0.36 0.117 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.558 0.058 0.576 0.122 ;
      RECT 0.45 0.058 0.468 0.122 ;
      RECT 0.288 0.058 0.306 0.122 ;
      RECT 0.18 0.022 0.198 0.086 ;
      RECT 0.072 0.022 0.09 0.086 ;
    LAYER M2 ;
      RECT 0.283 0.063 0.581 0.081 ;
      RECT 0.067 0.063 0.203 0.081 ;
    LAYER V1 ;
      RECT 0.558 0.063 0.576 0.081 ;
      RECT 0.45 0.063 0.468 0.081 ;
      RECT 0.288 0.063 0.306 0.081 ;
      RECT 0.18 0.063 0.198 0.081 ;
      RECT 0.072 0.063 0.09 0.081 ;
  END
END AOI22x1

MACRO BUFx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2 0 0 ;
  SIZE 0.27 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Y
END BUFx2

MACRO BUFx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END Y
END BUFx3

MACRO BUFx4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4 0 0 ;
  SIZE 0.378 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END Y
END BUFx4

MACRO BUFx8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8 0 0 ;
  SIZE 0.648 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END Y
END BUFx8

MACRO DFFHQNx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx1 0 0 ;
  SIZE 0.81 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.666 0.022 0.684 0.122 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END QN
  OBS
    LAYER M1 ;
      RECT 0.612 0.022 0.63 0.086 ;
      RECT 0.558 0.058 0.576 0.122 ;
      RECT 0.396 0.022 0.414 0.086 ;
    LAYER M2 ;
      RECT 0.391 0.063 0.581 0.081 ;
    LAYER V1 ;
      RECT 0.558 0.063 0.576 0.081 ;
      RECT 0.396 0.063 0.414 0.081 ;
  END
END DFFHQNx1

MACRO DFFHQNx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx2 0 0 ;
  SIZE 0.864 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.774 0.022 0.792 0.122 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.022 0.576 0.122 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END QN
  OBS
    LAYER M1 ;
      RECT 0.666 0.058 0.684 0.122 ;
      RECT 0.612 0.022 0.63 0.086 ;
      RECT 0.504 0.022 0.522 0.086 ;
      RECT 0.342 0.058 0.36 0.122 ;
    LAYER M2 ;
      RECT 0.337 0.063 0.689 0.081 ;
      RECT 0.499 0.027 0.635 0.045 ;
    LAYER V1 ;
      RECT 0.666 0.063 0.684 0.081 ;
      RECT 0.612 0.027 0.63 0.045 ;
      RECT 0.504 0.027 0.522 0.045 ;
      RECT 0.342 0.063 0.36 0.081 ;
  END
END DFFHQNx2

MACRO DFFHQNx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx3 0 0 ;
  SIZE 0.918 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.774 0.022 0.792 0.122 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END QN
  OBS
    LAYER M1 ;
      RECT 0.72 0.058 0.738 0.122 ;
      RECT 0.666 0.058 0.684 0.122 ;
      RECT 0.504 0.058 0.522 0.122 ;
    LAYER M2 ;
      RECT 0.499 0.063 0.689 0.081 ;
    LAYER V1 ;
      RECT 0.666 0.063 0.684 0.081 ;
      RECT 0.504 0.063 0.522 0.081 ;
  END
END DFFHQNx3

MACRO DHLx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx1 0 0 ;
  SIZE 0.594 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Q
  OBS
    LAYER M1 ;
      RECT 0.342 0.022 0.36 0.086 ;
      RECT 0.234 0.022 0.252 0.086 ;
    LAYER M2 ;
      RECT 0.229 0.063 0.365 0.081 ;
    LAYER V1 ;
      RECT 0.342 0.063 0.36 0.081 ;
      RECT 0.234 0.063 0.252 0.081 ;
  END
END DHLx1

MACRO DHLx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx2 0 0 ;
  SIZE 0.648 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.022 0.36 0.122 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Q
  OBS
    LAYER M1 ;
      RECT 0.396 0.058 0.414 0.122 ;
      RECT 0.288 0.058 0.306 0.122 ;
    LAYER M2 ;
      RECT 0.283 0.063 0.419 0.081 ;
    LAYER V1 ;
      RECT 0.396 0.063 0.414 0.081 ;
      RECT 0.288 0.063 0.306 0.081 ;
  END
END DHLx2

MACRO DHLx3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx3 0 0 ;
  SIZE 0.702 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.558 0.022 0.576 0.122 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Q
  OBS
    LAYER M1 ;
      RECT 0.504 0.058 0.522 0.122 ;
  END
END DHLx3

MACRO FAx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FAx1 0 0 ;
  SIZE 0.756 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.121 0.063 0.414 0.081 ;
      LAYER M1 ;
        RECT 0.396 0.022 0.414 0.086 ;
        RECT 0.126 0.022 0.144 0.122 ;
      LAYER V1 ;
        RECT 0.126 0.063 0.144 0.081 ;
        RECT 0.396 0.063 0.414 0.081 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.45 0.063 0.689 0.081 ;
      LAYER M1 ;
        RECT 0.666 0.058 0.684 0.122 ;
        RECT 0.45 0.022 0.468 0.122 ;
      LAYER V1 ;
        RECT 0.45 0.063 0.468 0.081 ;
        RECT 0.666 0.063 0.684 0.081 ;
    END
  END B
  PIN CI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.067 0.099 0.306 0.117 ;
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
        RECT 0.072 0.058 0.09 0.122 ;
      LAYER V1 ;
        RECT 0.072 0.099 0.09 0.117 ;
        RECT 0.288 0.099 0.306 0.117 ;
    END
  END CI
  PIN CON
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.342 0.099 0.527 0.117 ;
      LAYER M1 ;
        RECT 0.504 0.022 0.522 0.122 ;
        RECT 0.342 0.058 0.36 0.122 ;
      LAYER V1 ;
        RECT 0.342 0.099 0.36 0.117 ;
        RECT 0.504 0.099 0.522 0.117 ;
    END
  END CON
  PIN SN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END SN
END FAx1

MACRO INVx1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1 0 0 ;
  SIZE 0.162 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Y
END INVx1

MACRO INVx2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2 0 0 ;
  SIZE 0.216 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Y
END INVx2

MACRO INVx4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END Y
END INVx4

MACRO INVx8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8 0 0 ;
  SIZE 0.54 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.022 0.468 0.122 ;
    END
  END Y
END INVx8

MACRO NAND2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.058 0.198 0.122 ;
  END
END NAND2x1

MACRO NAND2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2 0 0 ;
  SIZE 0.54 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.022 0.468 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.504 0.058 0.522 0.122 ;
  END
END NAND2x2

MACRO NAND3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1 0 0 ;
  SIZE 0.594 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.022 0.36 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.022 0.522 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.175 0.063 0.311 0.081 ;
      LAYER M1 ;
        RECT 0.288 0.058 0.306 0.122 ;
        RECT 0.18 0.022 0.198 0.122 ;
      LAYER V1 ;
        RECT 0.18 0.063 0.198 0.081 ;
        RECT 0.288 0.063 0.306 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.022 0.414 0.086 ;
      RECT 0.234 0.022 0.252 0.086 ;
      RECT 0.018 0.022 0.036 0.086 ;
    LAYER M2 ;
      RECT 0.229 0.027 0.419 0.045 ;
    LAYER V1 ;
      RECT 0.396 0.027 0.414 0.045 ;
      RECT 0.234 0.027 0.252 0.045 ;
  END
END NAND3x1

MACRO NAND3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2 0 0 ;
  SIZE 1.08 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.022 0.63 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.283 0.027 0.959 0.045 ;
      LAYER M1 ;
        RECT 0.936 0.022 0.954 0.086 ;
        RECT 0.666 0.022 0.684 0.086 ;
        RECT 0.288 0.022 0.306 0.122 ;
      LAYER V1 ;
        RECT 0.288 0.027 0.306 0.045 ;
        RECT 0.666 0.027 0.684 0.045 ;
        RECT 0.936 0.027 0.954 0.045 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.99 0.022 1.008 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.823 0.099 1.067 0.117 ;
      LAYER M1 ;
        RECT 1.044 0.022 1.062 0.122 ;
        RECT 0.882 0.058 0.9 0.122 ;
        RECT 0.828 0.058 0.846 0.122 ;
      LAYER V1 ;
        RECT 0.828 0.099 0.846 0.117 ;
        RECT 0.882 0.099 0.9 0.117 ;
        RECT 1.044 0.099 1.062 0.117 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.72 0.058 0.738 0.122 ;
      RECT 0.342 0.058 0.36 0.122 ;
    LAYER M2 ;
      RECT 0.337 0.099 0.743 0.117 ;
    LAYER V1 ;
      RECT 0.72 0.099 0.738 0.117 ;
      RECT 0.342 0.099 0.36 0.117 ;
  END
END NAND3x2

MACRO NOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END Y
END NOR2x1

MACRO NOR2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2 0 0 ;
  SIZE 0.54 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Y
END NOR2x2

MACRO NOR3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1 0 0 ;
  SIZE 0.594 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.022 0.414 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.175 0.099 0.365 0.117 ;
      LAYER M1 ;
        RECT 0.342 0.058 0.36 0.122 ;
        RECT 0.18 0.022 0.198 0.122 ;
      LAYER V1 ;
        RECT 0.18 0.099 0.198 0.117 ;
        RECT 0.342 0.099 0.36 0.117 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.072 0.022 0.09 0.086 ;
  END
END NOR3x1

MACRO NOR3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2 0 0 ;
  SIZE 1.08 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.99 0.022 1.008 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.283 0.099 0.905 0.117 ;
      LAYER M1 ;
        RECT 0.882 0.022 0.9 0.122 ;
        RECT 0.666 0.058 0.684 0.122 ;
        RECT 0.288 0.058 0.306 0.122 ;
      LAYER V1 ;
        RECT 0.288 0.099 0.306 0.117 ;
        RECT 0.666 0.099 0.684 0.117 ;
        RECT 0.882 0.099 0.9 0.117 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.022 0.63 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.774 0.063 0.959 0.081 ;
      LAYER M1 ;
        RECT 0.936 0.022 0.954 0.122 ;
        RECT 0.828 0.022 0.846 0.086 ;
        RECT 0.774 0.022 0.792 0.086 ;
      LAYER V1 ;
        RECT 0.774 0.063 0.792 0.081 ;
        RECT 0.828 0.063 0.846 0.081 ;
        RECT 0.936 0.063 0.954 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.72 0.022 0.738 0.086 ;
      RECT 0.234 0.022 0.252 0.086 ;
    LAYER M2 ;
      RECT 0.229 0.063 0.738 0.081 ;
    LAYER V1 ;
      RECT 0.72 0.063 0.738 0.081 ;
      RECT 0.234 0.063 0.252 0.081 ;
  END
END NOR3x2

MACRO OAI21x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21x1 0 0 ;
  SIZE 0.486 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.283 0.063 0.419 0.081 ;
      LAYER M1 ;
        RECT 0.396 0.022 0.414 0.086 ;
        RECT 0.288 0.022 0.306 0.122 ;
      LAYER V1 ;
        RECT 0.288 0.063 0.306 0.081 ;
        RECT 0.396 0.063 0.414 0.081 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.342 0.022 0.36 0.086 ;
      RECT 0.18 0.022 0.198 0.086 ;
      RECT 0.018 0.022 0.036 0.086 ;
    LAYER M2 ;
      RECT 0.013 0.027 0.365 0.045 ;
    LAYER V1 ;
      RECT 0.342 0.027 0.36 0.045 ;
      RECT 0.18 0.027 0.198 0.045 ;
      RECT 0.018 0.027 0.036 0.045 ;
  END
END OAI21x1

MACRO OAI22x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22x1 0 0 ;
  SIZE 0.648 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.022 0.414 0.122 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.022 0.522 0.122 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.283 0.099 0.581 0.117 ;
      LAYER M1 ;
        RECT 0.558 0.058 0.576 0.122 ;
        RECT 0.45 0.022 0.468 0.122 ;
        RECT 0.288 0.058 0.306 0.122 ;
      LAYER V1 ;
        RECT 0.288 0.099 0.306 0.117 ;
        RECT 0.45 0.099 0.468 0.117 ;
        RECT 0.558 0.099 0.576 0.117 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.342 0.022 0.36 0.086 ;
      RECT 0.18 0.022 0.198 0.086 ;
      RECT 0.072 0.058 0.09 0.122 ;
    LAYER M2 ;
      RECT 0.067 0.063 0.365 0.081 ;
    LAYER V1 ;
      RECT 0.342 0.063 0.36 0.081 ;
      RECT 0.18 0.063 0.198 0.081 ;
      RECT 0.072 0.063 0.09 0.081 ;
  END
END OAI22x1

MACRO OR2x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Y
END OR2x2

MACRO OR3x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1 0 0 ;
  SIZE 0.324 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Y
END OR3x1

MACRO OR3x2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2 0 0 ;
  SIZE 0.378 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END Y
END OR3x2

MACRO XNOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x1 0 0 ;
  SIZE 0.594 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.022 0.522 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.121 0.063 0.473 0.081 ;
      LAYER M1 ;
        RECT 0.45 0.022 0.468 0.122 ;
        RECT 0.288 0.058 0.306 0.122 ;
        RECT 0.126 0.058 0.144 0.122 ;
      LAYER V1 ;
        RECT 0.126 0.063 0.144 0.081 ;
        RECT 0.288 0.063 0.306 0.081 ;
        RECT 0.45 0.063 0.468 0.081 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.558 0.022 0.576 0.086 ;
      RECT 0.396 0.022 0.414 0.086 ;
      RECT 0.342 0.058 0.36 0.122 ;
      RECT 0.234 0.022 0.252 0.086 ;
      RECT 0.072 0.058 0.09 0.122 ;
    LAYER M2 ;
      RECT 0.229 0.027 0.419 0.045 ;
      RECT 0.067 0.099 0.365 0.117 ;
    LAYER V1 ;
      RECT 0.396 0.027 0.414 0.045 ;
      RECT 0.342 0.099 0.36 0.117 ;
      RECT 0.234 0.027 0.252 0.045 ;
      RECT 0.072 0.099 0.09 0.117 ;
  END
END XNOR2x1

MACRO XOR2x1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x1 0 0 ;
  SIZE 0.594 BY 0.144 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.022 0.36 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.229 0.099 0.419 0.117 ;
      LAYER M1 ;
        RECT 0.396 0.058 0.414 0.122 ;
        RECT 0.234 0.022 0.252 0.122 ;
      LAYER V1 ;
        RECT 0.234 0.099 0.252 0.117 ;
        RECT 0.396 0.099 0.414 0.117 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 0.175 0.027 0.311 0.045 ;
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
        RECT 0.18 0.022 0.198 0.086 ;
      LAYER V1 ;
        RECT 0.18 0.027 0.198 0.045 ;
        RECT 0.288 0.027 0.306 0.045 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.45 0.022 0.468 0.086 ;
      RECT 0.126 0.058 0.144 0.122 ;
    LAYER M2 ;
      RECT 0.121 0.063 0.473 0.081 ;
    LAYER V1 ;
      RECT 0.45 0.063 0.468 0.081 ;
      RECT 0.126 0.063 0.144 0.081 ;
  END
END XOR2x1

END LIBRARY
