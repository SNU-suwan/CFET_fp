VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO AND2x2_ASAP7_75t_R_w4_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND2x2_ASAP7_75t_R_w4_8 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.058 0.252 0.158 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.058 0.144 0.158 ;
    END
  END Y
END AND2x2_ASAP7_75t_R_w4_8

MACRO AND3x1_ASAP7_75t_R_w4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x1_ASAP7_75t_R_w4_1 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.058 0.252 0.158 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.058 0.198 0.158 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END Y
END AND3x1_ASAP7_75t_R_w4_1

MACRO AND3x2_ASAP7_75t_R_w5_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AND3x2_ASAP7_75t_R_w5_0 0 0 ;
  SIZE 0.378 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.058 0.306 0.158 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END Y
END AND3x2_ASAP7_75t_R_w5_0

MACRO AOI21x1_ASAP7_75t_R_w6_3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI21x1_ASAP7_75t_R_w6_3 0 0 ;
  SIZE 0.27 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.238 0.09 0.338 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.202 0.198 0.302 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.126 0.022 0.144 0.338 ;
  END
END AOI21x1_ASAP7_75t_R_w6_3

MACRO AOI22x1_ASAP7_75t_R_w8_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22x1_ASAP7_75t_R_w8_0 0 0 ;
  SIZE 0.324 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.058 0.252 0.158 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.202 0.09 0.302 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.202 0.198 0.338 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.288 0.238 0.306 0.338 ;
      RECT 0.126 0.022 0.144 0.338 ;
  END
END AOI22x1_ASAP7_75t_R_w8_0

MACRO ASYNC_DFFHx1_ASAP7_75t_R_w22_19
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ASYNC_DFFHx1_ASAP7_75t_R_w22_19 0 0 ;
  SIZE 0.702 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.022 0.522 0.122 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.158 ;
    END
  END QN
  PIN RESET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.094 0.09 0.23 ;
    END
  END RESET
  PIN SET
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.612 0.022 0.63 0.122 ;
    END
  END SET
  OBS
    LAYER M1 ;
      RECT 0.612 0.202 0.63 0.302 ;
      RECT 0.558 0.022 0.576 0.086 ;
      RECT 0.558 0.13 0.576 0.338 ;
      RECT 0.504 0.202 0.522 0.302 ;
      RECT 0.45 0.022 0.468 0.23 ;
      RECT 0.45 0.274 0.468 0.338 ;
      RECT 0.396 0.058 0.414 0.266 ;
      RECT 0.342 0.022 0.36 0.338 ;
      RECT 0.288 0.022 0.306 0.086 ;
      RECT 0.288 0.13 0.306 0.302 ;
      RECT 0.234 0.022 0.252 0.086 ;
      RECT 0.234 0.13 0.252 0.23 ;
      RECT 0.234 0.274 0.252 0.338 ;
      RECT 0.18 0.202 0.198 0.266 ;
      RECT 0.126 0.058 0.144 0.338 ;
      RECT 0.072 0.274 0.09 0.338 ;
      RECT 0.018 0.274 0.036 0.338 ;
    LAYER M2 ;
      RECT 0.445 0.279 0.635 0.297 ;
      RECT 0.391 0.063 0.581 0.081 ;
      RECT 0.283 0.207 0.527 0.225 ;
      RECT 0.229 0.027 0.473 0.045 ;
      RECT 0.121 0.063 0.311 0.081 ;
      RECT 0.229 0.279 0.311 0.297 ;
      RECT 0.175 0.207 0.257 0.225 ;
      RECT 0.013 0.279 0.095 0.297 ;
    LAYER V1 ;
      RECT 0.612 0.279 0.63 0.297 ;
      RECT 0.558 0.063 0.576 0.081 ;
      RECT 0.504 0.207 0.522 0.225 ;
      RECT 0.45 0.027 0.468 0.045 ;
      RECT 0.45 0.279 0.468 0.297 ;
      RECT 0.396 0.063 0.414 0.081 ;
      RECT 0.288 0.063 0.306 0.081 ;
      RECT 0.288 0.207 0.306 0.225 ;
      RECT 0.288 0.279 0.306 0.297 ;
      RECT 0.234 0.027 0.252 0.045 ;
      RECT 0.234 0.207 0.252 0.225 ;
      RECT 0.234 0.279 0.252 0.297 ;
      RECT 0.18 0.207 0.198 0.225 ;
      RECT 0.126 0.063 0.144 0.081 ;
      RECT 0.072 0.279 0.09 0.297 ;
      RECT 0.018 0.279 0.036 0.297 ;
  END
END ASYNC_DFFHx1_ASAP7_75t_R_w22_19

MACRO BUFx2_ASAP7_75t_R_w3_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx2_ASAP7_75t_R_w3_0 0 0 ;
  SIZE 0.27 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.058 0.198 0.158 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Y
END BUFx2_ASAP7_75t_R_w3_0

MACRO BUFx3_ASAP7_75t_R_w4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx3_ASAP7_75t_R_w4_1 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.058 0.09 0.158 ;
    END
  END Y
END BUFx3_ASAP7_75t_R_w4_1

MACRO BUFx4_ASAP7_75t_R_w5_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx4_ASAP7_75t_R_w5_0 0 0 ;
  SIZE 0.378 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.058 0.198 0.158 ;
    END
  END Y
END BUFx4_ASAP7_75t_R_w5_0

MACRO BUFx8_ASAP7_75t_R_w10_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFx8_ASAP7_75t_R_w10_1 0 0 ;
  SIZE 0.648 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.058 0.144 0.158 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.022 0.414 0.122 ;
    END
  END Y
END BUFx8_ASAP7_75t_R_w10_1

MACRO DFFHQNx1_ASAP7_75t_R_w14_13
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx1_ASAP7_75t_R_w14_13 0 0 ;
  SIZE 0.486 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.094 0.414 0.23 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.022 0.36 0.122 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.238 0.036 0.338 ;
    END
  END QN
  OBS
    LAYER M1 ;
      RECT 0.234 0.13 0.252 0.338 ;
      RECT 0.18 0.022 0.198 0.23 ;
      RECT 0.126 0.058 0.144 0.266 ;
      RECT 0.072 0.094 0.09 0.23 ;
  END
END DFFHQNx1_ASAP7_75t_R_w14_13

MACRO DFFHQNx2_ASAP7_75t_R_w16_4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx2_ASAP7_75t_R_w16_4 0 0 ;
  SIZE 0.54 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.13 0.414 0.266 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.238 0.306 0.338 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.13 0.36 0.266 ;
    END
  END QN
  OBS
    LAYER M1 ;
      RECT 0.234 0.13 0.252 0.302 ;
      RECT 0.18 0.058 0.198 0.266 ;
      RECT 0.126 0.13 0.144 0.338 ;
      RECT 0.072 0.058 0.09 0.23 ;
  END
END DFFHQNx2_ASAP7_75t_R_w16_4

MACRO DFFHQNx3_ASAP7_75t_R_w16_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFFHQNx3_ASAP7_75t_R_w16_1 0 0 ;
  SIZE 0.54 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.238 0.144 0.338 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.202 0.468 0.302 ;
    END
  END D
  PIN QN
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.058 0.144 0.158 ;
    END
  END QN
  OBS
    LAYER M1 ;
      RECT 0.396 0.13 0.414 0.338 ;
      RECT 0.342 0.13 0.36 0.266 ;
      RECT 0.288 0.058 0.306 0.266 ;
      RECT 0.234 0.022 0.252 0.302 ;
      RECT 0.18 0.094 0.198 0.266 ;
  END
END DFFHQNx3_ASAP7_75t_R_w16_1

MACRO DHLx1_ASAP7_75t_R_w10_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DHLx1_ASAP7_75t_R_w10_1 0 0 ;
  SIZE 0.378 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.13 0.036 0.266 ;
    END
  END CLK
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.202 0.144 0.302 ;
    END
  END D
  PIN Q
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Q
  OBS
    LAYER M1 ;
      RECT 0.288 0.094 0.306 0.23 ;
      RECT 0.234 0.13 0.252 0.266 ;
      RECT 0.18 0.094 0.198 0.23 ;
      RECT 0.072 0.13 0.09 0.338 ;
  END
END DHLx1_ASAP7_75t_R_w10_1

MACRO INVx1_ASAP7_75t_R_w1_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx1_ASAP7_75t_R_w1_0 0 0 ;
  SIZE 0.162 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.158 ;
    END
  END Y
END INVx1_ASAP7_75t_R_w1_0

MACRO INVx2_ASAP7_75t_R_w2_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx2_ASAP7_75t_R_w2_1 0 0 ;
  SIZE 0.216 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.158 ;
    END
  END Y
END INVx2_ASAP7_75t_R_w2_1

MACRO INVx4_ASAP7_75t_R_w4_7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx4_ASAP7_75t_R_w4_7 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.058 0.252 0.158 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Y
END INVx4_ASAP7_75t_R_w4_7

MACRO INVx8_ASAP7_75t_R_w8_7
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVx8_ASAP7_75t_R_w8_7 0 0 ;
  SIZE 0.54 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.45 0.022 0.468 0.122 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.158 ;
    END
  END Y
END INVx8_ASAP7_75t_R_w8_7

MACRO NAND2x1_ASAP7_75t_R_w4_9
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x1_ASAP7_75t_R_w4_9 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.058 0.252 0.158 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END Y
END NAND2x1_ASAP7_75t_R_w4_9

MACRO NAND2x2_ASAP7_75t_R_w8_3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2x2_ASAP7_75t_R_w8_3 0 0 ;
  SIZE 0.324 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.238 0.144 0.338 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.18 0.094 0.198 0.23 ;
  END
END NAND2x2_ASAP7_75t_R_w8_3

MACRO NAND3x1_ASAP7_75t_R_w9_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x1_ASAP7_75t_R_w9_0 0 0 ;
  SIZE 0.594 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.058 0.36 0.158 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.058 0.522 0.158 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.022 0.414 0.122 ;
    END
  END Y
END NAND3x1_ASAP7_75t_R_w9_0

MACRO NAND3x2_ASAP7_75t_R_w18_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND3x2_ASAP7_75t_R_w18_0 0 0 ;
  SIZE 0.594 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.022 0.36 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.058 0.522 0.158 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.238 0.198 0.338 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.13 0.414 0.266 ;
      RECT 0.234 0.094 0.252 0.23 ;
  END
END NAND3x2_ASAP7_75t_R_w18_0

MACRO NOR2x1_ASAP7_75t_R_w4_9
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x1_ASAP7_75t_R_w4_9 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.158 ;
    END
  END Y
END NOR2x1_ASAP7_75t_R_w4_9

MACRO NOR2x2_ASAP7_75t_R_w8_3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2x2_ASAP7_75t_R_w8_3 0 0 ;
  SIZE 0.324 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.094 0.036 0.23 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.13 0.198 0.338 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.234 0.13 0.252 0.266 ;
      RECT 0.126 0.13 0.144 0.266 ;
  END
END NOR2x2_ASAP7_75t_R_w8_3

MACRO NOR3x1_ASAP7_75t_R_w9_3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x1_ASAP7_75t_R_w9_3 0 0 ;
  SIZE 0.594 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.058 0.522 0.158 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.058 0.36 0.158 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.058 0.09 0.158 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.022 0.144 0.122 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.45 0.022 0.468 0.158 ;
  END
END NOR3x1_ASAP7_75t_R_w9_3

MACRO NOR3x2_ASAP7_75t_R_w18_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR3x2_ASAP7_75t_R_w18_0 0 0 ;
  SIZE 0.594 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.094 0.522 0.23 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.342 0.238 0.36 0.338 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.13 0.198 0.266 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.202 0.09 0.302 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.396 0.094 0.414 0.338 ;
      RECT 0.234 0.13 0.252 0.338 ;
  END
END NOR3x2_ASAP7_75t_R_w18_0

MACRO OAI21x1_ASAP7_75t_R_w6_3
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI21x1_ASAP7_75t_R_w6_3 0 0 ;
  SIZE 0.27 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.13 0.198 0.266 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A2
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.238 0.09 0.338 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.202 0.036 0.302 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.126 0.13 0.144 0.302 ;
  END
END OAI21x1_ASAP7_75t_R_w6_3

MACRO OAI22x1_ASAP7_75t_R_w8_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22x1_ASAP7_75t_R_w8_0 0 0 ;
  SIZE 0.324 BY 0.36 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.238 0.09 0.338 ;
    END
  END A1
  PIN A2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.022 0.09 0.122 ;
    END
  END A2
  PIN B1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.238 0.198 0.338 ;
    END
  END B1
  PIN B2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END B2
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.094 0.036 0.23 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.234 0.022 0.252 0.338 ;
      RECT 0.126 0.13 0.144 0.302 ;
  END
END OAI22x1_ASAP7_75t_R_w8_0

MACRO OR2x2_ASAP7_75t_R_w4_8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR2x2_ASAP7_75t_R_w4_8 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.022 0.252 0.122 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.058 0.144 0.158 ;
    END
  END Y
END OR2x2_ASAP7_75t_R_w4_8

MACRO OR3x1_ASAP7_75t_R_w4_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x1_ASAP7_75t_R_w4_1 0 0 ;
  SIZE 0.324 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.058 0.252 0.158 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.022 0.198 0.122 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.126 0.058 0.144 0.158 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.158 ;
    END
  END Y
END OR3x1_ASAP7_75t_R_w4_1

MACRO OR3x2_ASAP7_75t_R_w5_0
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OR3x2_ASAP7_75t_R_w5_0 0 0 ;
  SIZE 0.378 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.288 0.022 0.306 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.234 0.058 0.252 0.158 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.058 0.198 0.158 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.072 0.058 0.09 0.158 ;
    END
  END Y
END OR3x2_ASAP7_75t_R_w5_0

MACRO XNOR2x1_ASAP7_75t_R_w9_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XNOR2x1_ASAP7_75t_R_w9_1 0 0 ;
  SIZE 0.594 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.504 0.022 0.522 0.122 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.058 0.198 0.158 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.022 0.036 0.122 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.45 0.022 0.468 0.086 ;
      RECT 0.342 0.022 0.36 0.086 ;
      RECT 0.288 0.058 0.306 0.122 ;
      RECT 0.126 0.022 0.144 0.086 ;
    LAYER M2 ;
      RECT 0.121 0.027 0.473 0.045 ;
      RECT 0.283 0.063 0.365 0.081 ;
    LAYER V1 ;
      RECT 0.45 0.027 0.468 0.045 ;
      RECT 0.342 0.063 0.36 0.081 ;
      RECT 0.288 0.063 0.306 0.081 ;
      RECT 0.126 0.027 0.144 0.045 ;
  END
END XNOR2x1_ASAP7_75t_R_w9_1

MACRO XOR2x1_ASAP7_75t_R_w9_1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR2x1_ASAP7_75t_R_w9_1 0 0 ;
  SIZE 0.594 BY 0.18 ;
  SYMMETRY X Y ;
  SITE coreSite ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.396 0.058 0.414 0.158 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.18 0.058 0.198 0.158 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 0.018 0.058 0.036 0.158 ;
    END
  END Y
  OBS
    LAYER M1 ;
      RECT 0.342 0.094 0.36 0.158 ;
      RECT 0.126 0.094 0.144 0.158 ;
    LAYER M2 ;
      RECT 0.121 0.135 0.365 0.153 ;
    LAYER V1 ;
      RECT 0.342 0.135 0.36 0.153 ;
      RECT 0.126 0.135 0.144 0.153 ;
  END
END XOR2x1_ASAP7_75t_R_w9_1

END LIBRARY
